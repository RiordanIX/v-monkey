module main

import (
	os
	repl
)

fn main() {
	println("Hello, this is the Monkey programming language!")
	repl.start()
}
